module BCD_counter (clk, reset, value);
	input clk, reset;
	output [19:0] value; //5 Digits
	
endmodule
