module BCD_counter #(parameter SIZE = 1)(clk, enable, value)

endmodule
