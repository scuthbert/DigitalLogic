module top(SW);
	input[9:0] SW;


endmodule
